module ddr3 (
    input wire clk,
    input wire rst,
    input wire [15:0] addr��
    input wire [1:0] ba
);
    
endmodule