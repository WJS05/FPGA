module ddr3 (
    input wire clk,
    input wire rst
);
    
endmodule